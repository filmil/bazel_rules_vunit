library vunit;

entity tb is
end entity;

architecture sim of tb is
begin
end architecture;
